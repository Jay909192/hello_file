module mux();
endmodule 

