module verilog 

input clk;
input rst;
endmodule 
