module verilog 
this is new feature;
input clk;
input rst;
endmodule
hello 

