module verilog 

input clk;
input rst;
input sequence_in;
output data_out;

endmodule 
