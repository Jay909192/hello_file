module adder ();
endmodule 
