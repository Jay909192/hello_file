module verilog( 
input clk,
input rst,
input sequence_in,
output data_out
);
always @( posedge clk or negedge rst)
begin
 
end

endmodule 
